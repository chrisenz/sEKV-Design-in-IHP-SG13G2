Simulation of the Miller OTA designed with the sEKV model

.lib /Simulations/models/cornerMOSlv.lib mos_tt ; model file for PSP
.include size_bias.par ; Size and bias values
.include pulse.par ; Pulse parameters for transient simulation
.include Miller_OTA.net ; Circuit netlist

.control
 op
 save v(out)
 write $inputdir/Miller_OTA.ac.op
* reset all
 ac dec 41 10 100MEG
 let AclmagdB=vdb(out)
 let Aclphdeg=180/PI*vp(out)
 let Aol=v(out)/(1-v(out))
 let AolmagdB=vdb(Aol)
 let Aolphdeg=180/PI*vp(Aol)
 meas ac fc when Aphdeg=-45
 set numdgt=12
 set wr_singlescale
 set wr_vecnames
* wrdata $inputdir/Miller_OTA.ac.dat AmagdB Aphdeg
 wrdata $inputdir/Miller_OTA.ac.dat vr(out) vi(out) AclmagdB Aclphdeg AolmagdB Aolphdeg
.endc
.end
