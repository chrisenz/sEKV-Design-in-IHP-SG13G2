OSDI PSP nMOS noise analysis

.lib /Simulations/models/cornerMOSlv.lib mos_tt
.include noise.par ; Size and bias values
.include noise.net ; Circuit netlist

.control
 op
 noise V(out) Vin dec $&decPts $&fmin $&fmax
 setplot noise1
 set wr_singlescale
 set wr_vecnames
 wrdata $inputdir/noise.dat inoise_spectrum onoise_spectrum
.endc
.end
