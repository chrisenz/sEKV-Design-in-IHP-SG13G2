Simulation of the symmetrical OTA designed with the sEKV model

.lib /Simulations/models/cornerMOSlv.lib mos_tt ; model file for PSP
.include size_bias.par ; Size and bias values
.include Miller_OTA.net ; Circuit netlist

.control
 op
 save v(out)
 write $inputdir/Miller_OTA.ac.op
* reset all
 ac dec 41 10 100MEG
 let AmagdB=vdb(out)
 let Aphdeg=180/PI*vp(out)
 meas ac Adc max AmagdB
 meas ac GBW when AmagdB=0
 meas ac PGBW find Aphdeg at=GBW
 set wr_singlescale
 set wr_vecnames
 wrdata $inputdir/Miller_OTA.ac.dat AmagdB Aphdeg
.endc
.end
