OSDI PSP nMOS noise analysis

.lib /Simulations/models/cornerMOSlv.lib mos_tt
.include noise.op.par ; Size and bias values
.include noise.net ; Circuit netlist

.control
 save @n.xp.Nsg13_lv_pmos[weff] @n.xp.Nsg13_lv_pmos[weff] @n.xp.Nsg13_lv_pmos[leff] @n.xp.Nsg13_lv_pmos[ids] @n.xp.Nsg13_lv_pmos[gm] @n.xp.Nsg13_lv_pmos[gds] @n.xp.Nsg13_lv_pmos[sid] @n.xp.Nsg13_lv_pmos[sqrtsfw] @n.xp.Nsg13_lv_pmos[sfl] @n.xp.Nsg13_lv_pmos[sqrtsff] @n.xp.Nsg13_lv_pmos[fknee]
 op
 wrnodev $inputdir/noise.op.ic
 set wr_singlescale
 set wr_vecnames
 wrdata $inputdir/noise.op.dat @n.xp.Nsg13_lv_pmos[weff] @n.xp.Nsg13_lv_pmos[leff] @n.xp.Nsg13_lv_pmos[ids] @n.xp.Nsg13_lv_pmos[gm] @n.xp.Nsg13_lv_pmos[gds] @n.xp.Nsg13_lv_pmos[sid] @n.xp.Nsg13_lv_pmos[sqrtsfw] @n.xp.Nsg13_lv_pmos[sfl] @n.xp.Nsg13_lv_pmos[sqrtsff] @n.xp.Nsg13_lv_pmos[fknee]
.endc
.end
