OSDI PSP nMOS VP-VG characteristic

.lib cornerMOSlv.lib mos_tt
.include vpvg.par ; Size and bias values
.include vpvg.net ; Circuit netlist

.control
 options GMIN=1e-15
 dc VG $&VGmin $&VGmax $&dVG
 let VP = v(s)
 meas dc VT0 WHEN V(s)=0.0
 set wr_singlescale
 set wr_vecnames
 wrdata $inputdir/vpvg.dat VP
.endc
.end
